rgb 0 0 0
s 0.5 0.5
M -49.49854 10.250898
l 0 -15.2894224
l 70.217363 0
L -10.425973 -27.972434
L 63.755273 2.6064096
L -10.425973 33.184808
l 31.144796 -22.93391
l -70.217363 0
f
