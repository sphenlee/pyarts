s 1 -1
rgb 0 0 0
M -4.2731748 -9.9571068
l -7.2985242 0
l 0 21.9999998
l 22.875 0
l 0 -21.9999998
l -8.1250001 0
l -7.4711941 0
l 0 7.8392046
l 7.7400388 0
l 0 -7.8223688
k

M -1.53125 -8.8281251
l 1.78125 0
l 0 5.546875
l -1.796875 0
l 0.015625 -5.546875
k

M -0.3125 0.06249998
C 0.85073904 0.10952916 1.9806289 0.70035869 2.6829458 1.6288455
C 3.3852627 2.5573323 3.6463073 3.8053652 3.375 4.9375
C 3.1812067 5.7461777 2.7244863 6.4900948 2.0890625 7.02652
C 1.4536387 7.5629453 0.64263413 7.8885845 -0.1875 7.9375
C -1.2404235 7.9995434 -2.311545 7.6077037 -3.079198 6.8843737
C -3.8468511 6.1610438 -4.3012718 5.1171901 -4.3125 4.0625
C -4.3236805 3.0122889 -3.8960804 1.9642266 -3.1534269 1.2215731
C -2.4107734 0.47891961 -1.3627111 0.05131944 -0.3125 0.06249998
k
