rgb 0 0 0
s 0.7 0.7
M 2.126468 10.792902
l 0 3.508804
l 12.373773 0
l 0 -11.944865
l -3.58346 0
l 0 8.436061
l -8.790313 0
f
M 2.232046 -10.99431
l 0 -3.508804
l 12.373773 0
l 0 11.9448647
l -3.583459 0
l 0 -8.4360607
l -8.790314 0
f
M -10.676801 -2.0006652
l -3.508804 0
l 0.05279 -12.3737728
l 11.9448651 0
l 0 3.58346
l -8.4360611 0
l -0.05279 8.7903128
f
M -1.894313 10.687324
l 0 3.508804
l -12.373773 0
l 0 -11.944865
l 3.58346 0
l 0 8.43606
l 8.790313 0
f
