rgb 0 0 0
s 0.5 0.5
M -22.394986 4.0998216
l 0 -7.4593421
L 15.007543 -3.633013
L 14.854824 -14.548424
L 32.858825 0.37025994
L 14.854824 15.288725
L 15.007543 3.8263292
l -37.402529 0.2734924
f