rgb 0 0 0
s 0.5 0.5
M -22.394986 4.0998216
l 0 -7.4593421
L 15.007543 -3.633013
L 14.854824 -14.548424
L 32.858825 0.37025994
L 14.854824 15.288725
L 15.007543 3.8263292
l -37.402529 0.2734924
f
M 20.0625 -23.75
C 6.880679 -23.75   -3.875 -12.994321   -3.875 0.1875
c 0 13.181821       10.755679 23.9375   23.9375 23.9375
C 33.244321 24.125  44 13.369321        44 0.1875
C 44 -12.994321     33.244321 -23.75    20.0625 -23.75
z
m 0 6.5
C 29.731461 -17.25  37.5 -9.4814605     37.5 0.1875
C 37.5 9.856461     29.731461 17.625    20.0625 17.625
C 10.393539 17.625  2.625 9.856461      2.625 0.1875
c 0 -9.6689605      7.768539 -17.4375   17.4375 -17.4375
z
f
