rgb 0 0 0
M 0.37880719 -9.5425235
L -5.555839 3.8419977
L 8.270624 10.155451
z
k